module stage1_64_tb #(
    parameter   WIDTH = 16
);
    reg clk;
    reg signed [(WIDTH*64)-1:0] x0_re, x0_im;
    wire signed [(WIDTH*64)-1:0] x1_re, x1_im;

    Stage1_64 dut (
        .x0_re(x0_re),
        .x0_im(x0_im),
        .x1_re(x1_re),
        .x1_im(x1_im)
    );

    always begin
        clk = 1'b0;
        forever #10 clk = ~clk;
    end

    initial begin
        x0_re = 64'b0;
        x0_im = 64'b0;

        #20

        x0_re = {
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000
        };

        x0_im = {
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000000000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000,
            16'b0000100000000000
        };
    end

endmodule